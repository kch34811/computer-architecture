module ALUControlUnit (input all_of_inst, output reg [2:0] alu_op);

    always @(all_of_inst) begin
        



    end

endmodule