module branch_predictor(input reset, 
                        input clk, 
                        input is_branch,
                        input [31:0] current_pc, 
                        input [31:0] next_pc,
                        );

  

endmodule